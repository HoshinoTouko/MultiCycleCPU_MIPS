library verilog;
use verilog.vl_types.all;
entity run is
end run;
